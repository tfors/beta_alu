`timescale 1ns/100ps

module alu_bool_tb;

reg clock = 0;

reg   [3:0] bfn;
reg  [31:0] a;
reg  [31:0] b;
wire [31:0] y;

// -------------------------------------------------------
// CLOCK GENERATION
// -------------------------------------------------------

always begin
	clock=0; #4;  // 125 MHz
	clock=1; #4;
end

// -------------------------------------------------------
// INITIALIZATION
// -------------------------------------------------------

initial begin
	if ($test$plusargs("vcd")) begin
		$dumpfile ("alu_bool_tb.vcd");
		$dumpvars (5, alu_bool_tb, dut);
	end
end

// -------------------------------------------------------
// TEST CASES
// -------------------------------------------------------

task test_case;
    input [67:0] inputs;
    input [31:0] expected_output;
    begin
        {bfn, a, b} <= inputs;
        @(posedge clock)
        if (y == expected_output) begin
            $display("pass: bfn=%01x, a=%08x, b=%08x => y=%08x",
                     inputs[67:64], inputs[63:32], inputs[31:0],
                     y);
        end else begin
            $error("FAIL: bfn=%01x, a=%08x, b=%08x => y=%08x (expected %08x)",
                   inputs[67:64], inputs[63:32], inputs[31:0],
                   y,
                   expected_output);
        end
    end
endtask

initial begin
    @(posedge clock);
    $display("");
    test_case({4'b0000, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, 32'b00000000000000000000000000000000); //  1: bfn=0b0000, a=0XFF00FF00, b=0XFFFF0000, y=0X00000000
    test_case({4'b0001, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, 32'b00000000000000000000000011111111); //  2: bfn=0b0001, a=0XFF00FF00, b=0XFFFF0000, y=0X000000FF
    test_case({4'b0010, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, 32'b00000000000000001111111100000000); //  3: bfn=0b0010, a=0XFF00FF00, b=0XFFFF0000, y=0X0000FF00
    test_case({4'b0011, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, 32'b00000000000000001111111111111111); //  4: bfn=0b0011, a=0XFF00FF00, b=0XFFFF0000, y=0X0000FFFF
    test_case({4'b0100, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, 32'b00000000111111110000000000000000); //  5: bfn=0b0100, a=0XFF00FF00, b=0XFFFF0000, y=0X00FF0000
    test_case({4'b0101, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, 32'b00000000111111110000000011111111); //  6: bfn=0b0101, a=0XFF00FF00, b=0XFFFF0000, y=0X00FF00FF
    test_case({4'b0110, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, 32'b00000000111111111111111100000000); //  7: bfn=0b0110, a=0XFF00FF00, b=0XFFFF0000, y=0X00FFFF00
    test_case({4'b0111, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, 32'b00000000111111111111111111111111); //  8: bfn=0b0111, a=0XFF00FF00, b=0XFFFF0000, y=0X00FFFFFF
    test_case({4'b1000, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, 32'b11111111000000000000000000000000); //  9: bfn=0b1000, a=0XFF00FF00, b=0XFFFF0000, y=0XFF000000
    test_case({4'b1001, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, 32'b11111111000000000000000011111111); // 10: bfn=0b1001, a=0XFF00FF00, b=0XFFFF0000, y=0XFF0000FF
    test_case({4'b1010, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, 32'b11111111000000001111111100000000); // 11: bfn=0b1010, a=0XFF00FF00, b=0XFFFF0000, y=0XFF00FF00
    test_case({4'b1011, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, 32'b11111111000000001111111111111111); // 12: bfn=0b1011, a=0XFF00FF00, b=0XFFFF0000, y=0XFF00FFFF
    test_case({4'b1100, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, 32'b11111111111111110000000000000000); // 13: bfn=0b1100, a=0XFF00FF00, b=0XFFFF0000, y=0XFFFF0000
    test_case({4'b1101, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, 32'b11111111111111110000000011111111); // 14: bfn=0b1101, a=0XFF00FF00, b=0XFFFF0000, y=0XFFFF00FF
    test_case({4'b1110, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, 32'b11111111111111111111111100000000); // 15: bfn=0b1110, a=0XFF00FF00, b=0XFFFF0000, y=0XFFFFFF00
    test_case({4'b1111, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, 32'b11111111111111111111111111111111); // 16: bfn=0b1111, a=0XFF00FF00, b=0XFFFF0000, y=0XFFFFFFFF
    $display("");
    $finish;
end


alu_bool dut (
    .bfn(bfn),
    .a(a),
    .b(b),
    .y(y)
);

endmodule
