`timescale 1ns/100ps

module cla_add32_tb;

reg clock = 0;

reg [31:0] a;
reg [31:0] b;
reg ci;
wire g;
wire p;
wire [31:0] s;

// -------------------------------------------------------
// CLOCK GENERATION
// -------------------------------------------------------

always begin
	clock=0; #4;  // 125 MHz
	clock=1; #4;
end

// -------------------------------------------------------
// INITIALIZATION
// -------------------------------------------------------

initial begin
	if ($test$plusargs("vcd")) begin
		$dumpfile ("cla_add32_tb.vcd");
		$dumpvars (5, cla_add32_tb, dut);
	end
end

// -------------------------------------------------------
// TEST CASES
// -------------------------------------------------------

task test_case;
    input [64:0] inputs;
    input [31:0] expected_output;
    begin
        {a, b, ci} <= inputs;
        @(posedge clock)
        if (s == expected_output) begin
            $display("pass: a=%08x, b=%08x, cin=%d => s=%08x",
                     inputs[64:33], inputs[32:1], inputs[0],
                     s);
        end else begin
            $error("FAIL: a=%08x, b=%08x, cin=%d => s=%08x (expected %08x)",
                   inputs[64:33], inputs[32:1], inputs[0],
                   s,
                   expected_output);
        end
    end
endtask

initial begin
    @(posedge clock);
    $display("");
    test_case({32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 1'b0}, 32'b00000000000000000000000000000000);
    test_case({32'b00000000000000000000000000000001, 32'b00000000000000000000000000000000, 1'b0}, 32'b00000000000000000000000000000001);
    test_case({32'b00000000000000000000000000000000, 32'b00000000000000000000000000000001, 1'b0}, 32'b00000000000000000000000000000001);
    test_case({32'b00000000000000000000000000000001, 32'b00000000000000000000000000000001, 1'b0}, 32'b00000000000000000000000000000010);
    test_case({32'b00000000000000000000000000000010, 32'b00000000000000000000000000000010, 1'b0}, 32'b00000000000000000000000000000100);
    test_case({32'b11111111111111111111111111111110, 32'b00000000000000000000000000000001, 1'b0}, 32'b11111111111111111111111111111111);
    test_case({32'b11111111111111111111111111111111, 32'b00000000000000000000000000000001, 1'b0}, 32'b00000000000000000000000000000000);
    test_case({32'b11111111111111111111111111111111, 32'b00000000000000000000000000000000, 1'b1}, 32'b00000000000000000000000000000000);
    test_case({32'b11111111111111110000000000000000, 32'b00000000000000001111111111111111, 1'b0}, 32'b11111111111111111111111111111111);
    test_case({32'b11111111111111110000000000000001, 32'b00000000000000001111111111111111, 1'b0}, 32'b00000000000000000000000000000000);
    test_case({32'b11111111111111110000000000000000, 32'b00000000000000001111111111111111, 1'b1}, 32'b00000000000000000000000000000000);
    test_case({32'b11111111111111110000000000000001, 32'b00000000000000001111111111111111, 1'b1}, 32'b00000000000000000000000000000001);
    $display("");
    $finish;
end


cla_add32 dut (
    .a(a),
    .b(b),
    .ci(ci),
    .g(g),
    .p(p),
    .s(s)
);

endmodule
