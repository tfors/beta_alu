`timescale 1ns/100ps

module beta_alu_tb;

reg clock = 0;

reg  [31:0] a;
reg  [31:0] b;
reg   [5:0] fn;
wire [31:0] y;

// -------------------------------------------------------
// CLOCK GENERATION
// -------------------------------------------------------

always begin
	clock=0; #4;  // 125 MHz
	clock=1; #4;
end

// -------------------------------------------------------
// INITIALIZATION
// -------------------------------------------------------

initial begin
	if ($test$plusargs("vcd")) begin
		$dumpfile ("beta_alu_tb.vcd");
		$dumpvars (5, beta_alu_tb, dut);
	end
end

// -------------------------------------------------------
// TEST CASES
// -------------------------------------------------------

task test_case;
    input [69:0] inputs;
    input [34:0] expected_output;
    begin
        {fn, a, b} <= inputs;
        @(posedge clock)
        if ({y, dut.z, dut.v, dut.n} == expected_output) begin
            $display("pass: fn=%02x, a=%08x, b=%08x => y=%08x, zvn=%01x",
                     inputs[69:64], inputs[63:32], inputs[31:0],
                     y, {dut.z, dut.v, dut.n});
        end else begin
            $error("FAIL: fn=%02x, a=%08x, b=%02x => y=%08x, zvn=%01x (expected %08x, %01x)",
                   inputs[69:64], inputs[63:32], inputs[31:0],
                   y, {dut.z, dut.v, dut.n},
                   expected_output[34:3], expected_output[2:0]);
        end
    end
endtask

initial begin
	@(posedge clock);
	$display("");
	test_case({6'b100010, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b00000000000000001111111100000000, 3'b001}); //   3: fn=F0010, a=0xff00ff00, b=0xffff0000, y=0x0000ff00
	test_case({6'b100001, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b00000000000000000000000011111111, 3'b001}); //   2: fn=F0001, a=0xff00ff00, b=0xffff0000, y=0x000000ff
	test_case({6'b100011, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b00000000000000001111111111111111, 3'b001}); //   4: fn=F0011, a=0xff00ff00, b=0xffff0000, y=0x0000ffff
	test_case({6'b100100, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b00000000111111110000000000000000, 3'b001}); //   5: fn=F0100, a=0xff00ff00, b=0xffff0000, y=0x00ff0000
	test_case({6'b100101, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b00000000111111110000000011111111, 3'b001}); //   6: fn=F0101, a=0xff00ff00, b=0xffff0000, y=0x00ff00ff
	test_case({6'b100110, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b00000000111111111111111100000000, 3'b001}); //   7: fn=  XOR, a=0xff00ff00, b=0xffff0000, y=0x00ffff00
	test_case({6'b100111, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b00000000111111111111111111111111, 3'b001}); //   8: fn=F0111, a=0xff00ff00, b=0xffff0000, y=0x00ffffff
	test_case({6'b101000, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b11111111000000000000000000000000, 3'b001}); //   9: fn=  AND, a=0xff00ff00, b=0xffff0000, y=0xff000000
	test_case({6'b100000, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b00000000000000000000000000000000, 3'b001}); //   1: fn=F0000, a=0xff00ff00, b=0xffff0000, y=0x00000000
	test_case({6'b101001, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b11111111000000000000000011111111, 3'b001}); //  10: fn= XNOR, a=0xff00ff00, b=0xffff0000, y=0xff0000ff
	test_case({6'b101010, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b11111111000000001111111100000000, 3'b001}); //  11: fn=    A, a=0xff00ff00, b=0xffff0000, y=0xff00ff00
	test_case({6'b101011, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b11111111000000001111111111111111, 3'b001}); //  12: fn=F1011, a=0xff00ff00, b=0xffff0000, y=0xff00ffff
	test_case({6'b101100, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b11111111111111110000000000000000, 3'b001}); //  13: fn=F1100, a=0xff00ff00, b=0xffff0000, y=0xffff0000
	test_case({6'b101101, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b11111111111111110000000011111111, 3'b001}); //  14: fn=F1101, a=0xff00ff00, b=0xffff0000, y=0xffff00ff
	test_case({6'b101110, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b11111111111111111111111100000000, 3'b001}); //  15: fn=   OR, a=0xff00ff00, b=0xffff0000, y=0xffffff00
	test_case({6'b101111, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b11111111111111111111111111111111, 3'b001}); //  16: fn=F1111, a=0xff00ff00, b=0xffff0000, y=0xffffffff
	test_case({6'b110000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000000, 3'b100}); //  17: fn=  SHL, a=0x00000000, b=0x00000000, y=0x00000000
	test_case({6'b110001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000000, 3'b100}); //  18: fn=  SHR, a=0x00000000, b=0x00000000, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000000, 3'b100}); //  19: fn=  SRA, a=0x00000000, b=0x00000000, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000000, 3'b000}); //  20: fn=  SHL, a=0x00000000, b=0x00000001, y=0x00000000
	test_case({6'b110001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000000, 3'b001}); //  21: fn=  SHR, a=0x00000000, b=0x00000001, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000000, 3'b001}); //  22: fn=  SRA, a=0x00000000, b=0x00000001, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000010}, {32'b00000000000000000000000000000000, 3'b000}); //  23: fn=  SHL, a=0x00000000, b=0x00000002, y=0x00000000
	test_case({6'b110001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000010}, {32'b00000000000000000000000000000000, 3'b001}); //  24: fn=  SHR, a=0x00000000, b=0x00000002, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000010}, {32'b00000000000000000000000000000000, 3'b001}); //  25: fn=  SRA, a=0x00000000, b=0x00000002, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000100}, {32'b00000000000000000000000000000000, 3'b000}); //  26: fn=  SHL, a=0x00000000, b=0x00000004, y=0x00000000
	test_case({6'b110001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000100}, {32'b00000000000000000000000000000000, 3'b001}); //  27: fn=  SHR, a=0x00000000, b=0x00000004, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000100}, {32'b00000000000000000000000000000000, 3'b001}); //  28: fn=  SRA, a=0x00000000, b=0x00000004, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000001000}, {32'b00000000000000000000000000000000, 3'b000}); //  29: fn=  SHL, a=0x00000000, b=0x00000008, y=0x00000000
	test_case({6'b110001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000001000}, {32'b00000000000000000000000000000000, 3'b001}); //  30: fn=  SHR, a=0x00000000, b=0x00000008, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000001000}, {32'b00000000000000000000000000000000, 3'b001}); //  31: fn=  SRA, a=0x00000000, b=0x00000008, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000010000}, {32'b00000000000000000000000000000000, 3'b000}); //  32: fn=  SHL, a=0x00000000, b=0x00000010, y=0x00000000
	test_case({6'b110001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000010000}, {32'b00000000000000000000000000000000, 3'b001}); //  33: fn=  SHR, a=0x00000000, b=0x00000010, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000010000}, {32'b00000000000000000000000000000000, 3'b001}); //  34: fn=  SRA, a=0x00000000, b=0x00000010, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000000, 3'b000}); //  35: fn=  SHL, a=0x00000000, b=0x0000001f, y=0x00000000
	test_case({6'b110001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000000, 3'b001}); //  36: fn=  SHR, a=0x00000000, b=0x0000001f, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000000, 3'b001}); //  37: fn=  SRA, a=0x00000000, b=0x0000001f, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000001, 3'b000}); //  38: fn=  SHL, a=0x00000001, b=0x00000000, y=0x00000001
	test_case({6'b110001, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000001, 3'b000}); //  39: fn=  SHR, a=0x00000001, b=0x00000000, y=0x00000001
	test_case({6'b110011, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000001, 3'b000}); //  40: fn=  SRA, a=0x00000001, b=0x00000000, y=0x00000001
	test_case({6'b110000, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000010, 3'b000}); //  41: fn=  SHL, a=0x00000001, b=0x00000001, y=0x00000002
	test_case({6'b110001, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000000, 3'b100}); //  42: fn=  SHR, a=0x00000001, b=0x00000001, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000000, 3'b100}); //  43: fn=  SRA, a=0x00000001, b=0x00000001, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000010}, {32'b00000000000000000000000000000100, 3'b000}); //  44: fn=  SHL, a=0x00000001, b=0x00000002, y=0x00000004
	test_case({6'b110001, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000010}, {32'b00000000000000000000000000000000, 3'b001}); //  45: fn=  SHR, a=0x00000001, b=0x00000002, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000010}, {32'b00000000000000000000000000000000, 3'b001}); //  46: fn=  SRA, a=0x00000001, b=0x00000002, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000100}, {32'b00000000000000000000000000010000, 3'b000}); //  47: fn=  SHL, a=0x00000001, b=0x00000004, y=0x00000010
	test_case({6'b110001, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000100}, {32'b00000000000000000000000000000000, 3'b001}); //  48: fn=  SHR, a=0x00000001, b=0x00000004, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000100}, {32'b00000000000000000000000000000000, 3'b001}); //  49: fn=  SRA, a=0x00000001, b=0x00000004, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000001000}, {32'b00000000000000000000000100000000, 3'b000}); //  50: fn=  SHL, a=0x00000001, b=0x00000008, y=0x00000100
	test_case({6'b110001, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000001000}, {32'b00000000000000000000000000000000, 3'b001}); //  51: fn=  SHR, a=0x00000001, b=0x00000008, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000001000}, {32'b00000000000000000000000000000000, 3'b001}); //  52: fn=  SRA, a=0x00000001, b=0x00000008, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000010000}, {32'b00000000000000010000000000000000, 3'b000}); //  53: fn=  SHL, a=0x00000001, b=0x00000010, y=0x00010000
	test_case({6'b110001, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000010000}, {32'b00000000000000000000000000000000, 3'b001}); //  54: fn=  SHR, a=0x00000001, b=0x00000010, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000010000}, {32'b00000000000000000000000000000000, 3'b001}); //  55: fn=  SRA, a=0x00000001, b=0x00000010, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000011111}, {32'b10000000000000000000000000000000, 3'b000}); //  56: fn=  SHL, a=0x00000001, b=0x0000001f, y=0x80000000
	test_case({6'b110001, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000000, 3'b001}); //  57: fn=  SHR, a=0x00000001, b=0x0000001f, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000000, 3'b001}); //  58: fn=  SRA, a=0x00000001, b=0x0000001f, y=0x00000000
	test_case({6'b110000, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000000}, {32'b11111111111111111111111111111111, 3'b001}); //  59: fn=  SHL, a=0xffffffff, b=0x00000000, y=0xffffffff
	test_case({6'b110001, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000000}, {32'b11111111111111111111111111111111, 3'b001}); //  60: fn=  SHR, a=0xffffffff, b=0x00000000, y=0xffffffff
	test_case({6'b110011, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000000}, {32'b11111111111111111111111111111111, 3'b001}); //  61: fn=  SRA, a=0xffffffff, b=0x00000000, y=0xffffffff
	test_case({6'b110000, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000001}, {32'b11111111111111111111111111111110, 3'b100}); //  62: fn=  SHL, a=0xffffffff, b=0x00000001, y=0xfffffffe
	test_case({6'b110001, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000001}, {32'b01111111111111111111111111111111, 3'b001}); //  63: fn=  SHR, a=0xffffffff, b=0x00000001, y=0x7fffffff
	test_case({6'b110011, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000001}, {32'b11111111111111111111111111111111, 3'b001}); //  64: fn=  SRA, a=0xffffffff, b=0x00000001, y=0xffffffff
	test_case({6'b110000, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000010}, {32'b11111111111111111111111111111100, 3'b000}); //  65: fn=  SHL, a=0xffffffff, b=0x00000002, y=0xfffffffc
	test_case({6'b110001, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000010}, {32'b00111111111111111111111111111111, 3'b001}); //  66: fn=  SHR, a=0xffffffff, b=0x00000002, y=0x3fffffff
	test_case({6'b110011, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000010}, {32'b11111111111111111111111111111111, 3'b001}); //  67: fn=  SRA, a=0xffffffff, b=0x00000002, y=0xffffffff
	test_case({6'b110000, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000100}, {32'b11111111111111111111111111110000, 3'b000}); //  68: fn=  SHL, a=0xffffffff, b=0x00000004, y=0xfffffff0
	test_case({6'b110001, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000100}, {32'b00001111111111111111111111111111, 3'b001}); //  69: fn=  SHR, a=0xffffffff, b=0x00000004, y=0x0fffffff
	test_case({6'b110011, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000100}, {32'b11111111111111111111111111111111, 3'b001}); //  70: fn=  SRA, a=0xffffffff, b=0x00000004, y=0xffffffff
	test_case({6'b110000, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000001000}, {32'b11111111111111111111111100000000, 3'b000}); //  71: fn=  SHL, a=0xffffffff, b=0x00000008, y=0xffffff00
	test_case({6'b110001, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000001000}, {32'b00000000111111111111111111111111, 3'b001}); //  72: fn=  SHR, a=0xffffffff, b=0x00000008, y=0x00ffffff
	test_case({6'b110011, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000001000}, {32'b11111111111111111111111111111111, 3'b001}); //  73: fn=  SRA, a=0xffffffff, b=0x00000008, y=0xffffffff
	test_case({6'b110000, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000010000}, {32'b11111111111111110000000000000000, 3'b000}); //  74: fn=  SHL, a=0xffffffff, b=0x00000010, y=0xffff0000
	test_case({6'b110001, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000010000}, {32'b00000000000000001111111111111111, 3'b001}); //  75: fn=  SHR, a=0xffffffff, b=0x00000010, y=0x0000ffff
	test_case({6'b110011, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000010000}, {32'b11111111111111111111111111111111, 3'b001}); //  76: fn=  SRA, a=0xffffffff, b=0x00000010, y=0xffffffff
	test_case({6'b110000, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000011111}, {32'b10000000000000000000000000000000, 3'b000}); //  77: fn=  SHL, a=0xffffffff, b=0x0000001f, y=0x80000000
	test_case({6'b110001, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000001, 3'b001}); //  78: fn=  SHR, a=0xffffffff, b=0x0000001f, y=0x00000001
	test_case({6'b110011, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000011111}, {32'b11111111111111111111111111111111, 3'b001}); //  79: fn=  SRA, a=0xffffffff, b=0x0000001f, y=0xffffffff
	test_case({6'b110000, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000000}, {32'b00010010001101000101011001111000, 3'b000}); //  80: fn=  SHL, a=0x12345678, b=0x00000000, y=0x12345678
	test_case({6'b110001, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000000}, {32'b00010010001101000101011001111000, 3'b000}); //  81: fn=  SHR, a=0x12345678, b=0x00000000, y=0x12345678
	test_case({6'b110011, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000000}, {32'b00010010001101000101011001111000, 3'b000}); //  82: fn=  SRA, a=0x12345678, b=0x00000000, y=0x12345678
	test_case({6'b110000, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000001}, {32'b00100100011010001010110011110000, 3'b000}); //  83: fn=  SHL, a=0x12345678, b=0x00000001, y=0x2468acf0
	test_case({6'b110001, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000001}, {32'b00001001000110100010101100111100, 3'b000}); //  84: fn=  SHR, a=0x12345678, b=0x00000001, y=0x091a2b3c
	test_case({6'b110011, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000001}, {32'b00001001000110100010101100111100, 3'b000}); //  85: fn=  SRA, a=0x12345678, b=0x00000001, y=0x091a2b3c
	test_case({6'b110000, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000010}, {32'b01001000110100010101100111100000, 3'b000}); //  86: fn=  SHL, a=0x12345678, b=0x00000002, y=0x48d159e0
	test_case({6'b110001, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000010}, {32'b00000100100011010001010110011110, 3'b000}); //  87: fn=  SHR, a=0x12345678, b=0x00000002, y=0x048d159e
	test_case({6'b110011, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000010}, {32'b00000100100011010001010110011110, 3'b000}); //  88: fn=  SRA, a=0x12345678, b=0x00000002, y=0x048d159e
	test_case({6'b110000, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000100}, {32'b00100011010001010110011110000000, 3'b000}); //  89: fn=  SHL, a=0x12345678, b=0x00000004, y=0x23456780
	test_case({6'b110001, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000100}, {32'b00000001001000110100010101100111, 3'b000}); //  90: fn=  SHR, a=0x12345678, b=0x00000004, y=0x01234567
	test_case({6'b110011, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000100}, {32'b00000001001000110100010101100111, 3'b000}); //  91: fn=  SRA, a=0x12345678, b=0x00000004, y=0x01234567
	test_case({6'b110000, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000001000}, {32'b00110100010101100111100000000000, 3'b000}); //  92: fn=  SHL, a=0x12345678, b=0x00000008, y=0x34567800
	test_case({6'b110001, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000001000}, {32'b00000000000100100011010001010110, 3'b000}); //  93: fn=  SHR, a=0x12345678, b=0x00000008, y=0x00123456
	test_case({6'b110011, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000001000}, {32'b00000000000100100011010001010110, 3'b000}); //  94: fn=  SRA, a=0x12345678, b=0x00000008, y=0x00123456
	test_case({6'b110000, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000010000}, {32'b01010110011110000000000000000000, 3'b000}); //  95: fn=  SHL, a=0x12345678, b=0x00000010, y=0x56780000
	test_case({6'b110001, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000010000}, {32'b00000000000000000001001000110100, 3'b000}); //  96: fn=  SHR, a=0x12345678, b=0x00000010, y=0x00001234
	test_case({6'b110011, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000010000}, {32'b00000000000000000001001000110100, 3'b000}); //  97: fn=  SRA, a=0x12345678, b=0x00000010, y=0x00001234
	test_case({6'b110000, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000000, 3'b000}); //  98: fn=  SHL, a=0x12345678, b=0x0000001f, y=0x00000000
	test_case({6'b110001, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000000, 3'b000}); //  99: fn=  SHR, a=0x12345678, b=0x0000001f, y=0x00000000
	test_case({6'b110011, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000000, 3'b000}); // 100: fn=  SRA, a=0x12345678, b=0x0000001f, y=0x00000000
	test_case({6'b110000, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000000}, {32'b11111110110111001010101110011000, 3'b001}); // 101: fn=  SHL, a=0xfedcab98, b=0x00000000, y=0xfedcab98
	test_case({6'b110001, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000000}, {32'b11111110110111001010101110011000, 3'b001}); // 102: fn=  SHR, a=0xfedcab98, b=0x00000000, y=0xfedcab98
	test_case({6'b110011, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000000}, {32'b11111110110111001010101110011000, 3'b001}); // 103: fn=  SRA, a=0xfedcab98, b=0x00000000, y=0xfedcab98
	test_case({6'b110000, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000001}, {32'b11111101101110010101011100110000, 3'b001}); // 104: fn=  SHL, a=0xfedcab98, b=0x00000001, y=0xfdb95730
	test_case({6'b110001, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000001}, {32'b01111111011011100101010111001100, 3'b001}); // 105: fn=  SHR, a=0xfedcab98, b=0x00000001, y=0x7f6e55cc
	test_case({6'b110011, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000001}, {32'b11111111011011100101010111001100, 3'b001}); // 106: fn=  SRA, a=0xfedcab98, b=0x00000001, y=0xff6e55cc
	test_case({6'b110000, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000010}, {32'b11111011011100101010111001100000, 3'b001}); // 107: fn=  SHL, a=0xfedcab98, b=0x00000002, y=0xfb72ae60
	test_case({6'b110001, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000010}, {32'b00111111101101110010101011100110, 3'b001}); // 108: fn=  SHR, a=0xfedcab98, b=0x00000002, y=0x3fb72ae6
	test_case({6'b110011, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000010}, {32'b11111111101101110010101011100110, 3'b001}); // 109: fn=  SRA, a=0xfedcab98, b=0x00000002, y=0xffb72ae6
	test_case({6'b110000, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000100}, {32'b11101101110010101011100110000000, 3'b001}); // 110: fn=  SHL, a=0xfedcab98, b=0x00000004, y=0xedcab980
	test_case({6'b110001, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000100}, {32'b00001111111011011100101010111001, 3'b001}); // 111: fn=  SHR, a=0xfedcab98, b=0x00000004, y=0x0fedcab9
	test_case({6'b110011, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000100}, {32'b11111111111011011100101010111001, 3'b001}); // 112: fn=  SRA, a=0xfedcab98, b=0x00000004, y=0xffedcab9
	test_case({6'b110000, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000001000}, {32'b11011100101010111001100000000000, 3'b001}); // 113: fn=  SHL, a=0xfedcab98, b=0x00000008, y=0xdcab9800
	test_case({6'b110001, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000001000}, {32'b00000000111111101101110010101011, 3'b001}); // 114: fn=  SHR, a=0xfedcab98, b=0x00000008, y=0x00fedcab
	test_case({6'b110011, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000001000}, {32'b11111111111111101101110010101011, 3'b001}); // 115: fn=  SRA, a=0xfedcab98, b=0x00000008, y=0xfffedcab
	test_case({6'b110000, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000010000}, {32'b10101011100110000000000000000000, 3'b001}); // 116: fn=  SHL, a=0xfedcab98, b=0x00000010, y=0xab980000
	test_case({6'b110001, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000010000}, {32'b00000000000000001111111011011100, 3'b001}); // 117: fn=  SHR, a=0xfedcab98, b=0x00000010, y=0x0000fedc
	test_case({6'b110011, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000010000}, {32'b11111111111111111111111011011100, 3'b001}); // 118: fn=  SRA, a=0xfedcab98, b=0x00000010, y=0xfffffedc
	test_case({6'b110000, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000000, 3'b001}); // 119: fn=  SHL, a=0xfedcab98, b=0x0000001f, y=0x00000000
	test_case({6'b110001, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000001, 3'b001}); // 120: fn=  SHR, a=0xfedcab98, b=0x0000001f, y=0x00000001
	test_case({6'b110011, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000011111}, {32'b11111111111111111111111111111111, 3'b001}); // 121: fn=  SRA, a=0xfedcab98, b=0x0000001f, y=0xffffffff
	test_case({6'b010000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000000, 3'b100}); // 122: fn=  ADD, a=0x00000000, b=0x00000000, y=0x00000000
	test_case({6'b010000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000001, 3'b000}); // 123: fn=  ADD, a=0x00000000, b=0x00000001, y=0x00000001
	test_case({6'b010000, 32'b00000000000000000000000000000000, 32'b11111111111111111111111111111111}, {32'b11111111111111111111111111111111, 3'b001}); // 124: fn=  ADD, a=0x00000000, b=0x-0000001, y=0xffffffff
	test_case({6'b010000, 32'b00000000000000000000000000000000, 32'b10101010101010101010101010101010}, {32'b10101010101010101010101010101010, 3'b001}); // 125: fn=  ADD, a=0x00000000, b=0xaaaaaaaa, y=0xaaaaaaaa
	test_case({6'b010000, 32'b00000000000000000000000000000000, 32'b01010101010101010101010101010101}, {32'b01010101010101010101010101010101, 3'b000}); // 126: fn=  ADD, a=0x00000000, b=0x55555555, y=0x55555555
	test_case({6'b010000, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000001, 3'b000}); // 127: fn=  ADD, a=0x00000001, b=0x00000000, y=0x00000001
	test_case({6'b010000, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000010, 3'b000}); // 128: fn=  ADD, a=0x00000001, b=0x00000001, y=0x00000002
	test_case({6'b010000, 32'b00000000000000000000000000000001, 32'b11111111111111111111111111111111}, {32'b00000000000000000000000000000000, 3'b100}); // 129: fn=  ADD, a=0x00000001, b=0x-0000001, y=0x00000000
	test_case({6'b010000, 32'b00000000000000000000000000000001, 32'b10101010101010101010101010101010}, {32'b10101010101010101010101010101011, 3'b001}); // 130: fn=  ADD, a=0x00000001, b=0xaaaaaaaa, y=0xaaaaaaab
	test_case({6'b010000, 32'b00000000000000000000000000000001, 32'b01010101010101010101010101010101}, {32'b01010101010101010101010101010110, 3'b000}); // 131: fn=  ADD, a=0x00000001, b=0x55555555, y=0x55555556
	test_case({6'b010000, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000000}, {32'b11111111111111111111111111111111, 3'b001}); // 132: fn=  ADD, a=0x-0000001, b=0x00000000, y=0xffffffff
	test_case({6'b010000, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000000, 3'b100}); // 133: fn=  ADD, a=0x-0000001, b=0x00000001, y=0x00000000
	test_case({6'b010000, 32'b11111111111111111111111111111111, 32'b11111111111111111111111111111111}, {32'b11111111111111111111111111111110, 3'b001}); // 134: fn=  ADD, a=0x-0000001, b=0x-0000001, y=0xfffffffe
	test_case({6'b010000, 32'b11111111111111111111111111111111, 32'b10101010101010101010101010101010}, {32'b10101010101010101010101010101001, 3'b001}); // 135: fn=  ADD, a=0x-0000001, b=0xaaaaaaaa, y=0xaaaaaaa9
	test_case({6'b010000, 32'b11111111111111111111111111111111, 32'b01010101010101010101010101010101}, {32'b01010101010101010101010101010100, 3'b000}); // 136: fn=  ADD, a=0x-0000001, b=0x55555555, y=0x55555554
	test_case({6'b010000, 32'b10101010101010101010101010101010, 32'b00000000000000000000000000000000}, {32'b10101010101010101010101010101010, 3'b001}); // 137: fn=  ADD, a=0xaaaaaaaa, b=0x00000000, y=0xaaaaaaaa
	test_case({6'b010000, 32'b10101010101010101010101010101010, 32'b00000000000000000000000000000001}, {32'b10101010101010101010101010101011, 3'b001}); // 138: fn=  ADD, a=0xaaaaaaaa, b=0x00000001, y=0xaaaaaaab
	test_case({6'b010000, 32'b10101010101010101010101010101010, 32'b11111111111111111111111111111111}, {32'b10101010101010101010101010101001, 3'b001}); // 139: fn=  ADD, a=0xaaaaaaaa, b=0x-0000001, y=0xaaaaaaa9
	test_case({6'b010000, 32'b10101010101010101010101010101010, 32'b10101010101010101010101010101010}, {32'b01010101010101010101010101010100, 3'b010}); // 140: fn=  ADD, a=0xaaaaaaaa, b=0xaaaaaaaa, y=0x55555554
	test_case({6'b010000, 32'b10101010101010101010101010101010, 32'b01010101010101010101010101010101}, {32'b11111111111111111111111111111111, 3'b001}); // 141: fn=  ADD, a=0xaaaaaaaa, b=0x55555555, y=0xffffffff
	test_case({6'b010000, 32'b01010101010101010101010101010101, 32'b00000000000000000000000000000000}, {32'b01010101010101010101010101010101, 3'b000}); // 142: fn=  ADD, a=0x55555555, b=0x00000000, y=0x55555555
	test_case({6'b010000, 32'b01010101010101010101010101010101, 32'b00000000000000000000000000000001}, {32'b01010101010101010101010101010110, 3'b000}); // 143: fn=  ADD, a=0x55555555, b=0x00000001, y=0x55555556
	test_case({6'b010000, 32'b01010101010101010101010101010101, 32'b11111111111111111111111111111111}, {32'b01010101010101010101010101010100, 3'b000}); // 144: fn=  ADD, a=0x55555555, b=0x-0000001, y=0x55555554
	test_case({6'b010000, 32'b01010101010101010101010101010101, 32'b10101010101010101010101010101010}, {32'b11111111111111111111111111111111, 3'b001}); // 145: fn=  ADD, a=0x55555555, b=0xaaaaaaaa, y=0xffffffff
	test_case({6'b010000, 32'b01010101010101010101010101010101, 32'b01010101010101010101010101010101}, {32'b10101010101010101010101010101010, 3'b011}); // 146: fn=  ADD, a=0x55555555, b=0x55555555, y=0xaaaaaaaa
	test_case({6'b010001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000000, 3'b100}); // 147: fn=  SUB, a=0x00000000, b=0x00000000, y=0x00000000
	test_case({6'b010001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000001}, {32'b11111111111111111111111111111111, 3'b001}); // 148: fn=  SUB, a=0x00000000, b=0x00000001, y=0xffffffff
	test_case({6'b010001, 32'b00000000000000000000000000000000, 32'b11111111111111111111111111111111}, {32'b00000000000000000000000000000001, 3'b000}); // 149: fn=  SUB, a=0x00000000, b=0x-0000001, y=0x00000001
	test_case({6'b010001, 32'b00000000000000000000000000000000, 32'b10101010101010101010101010101010}, {32'b01010101010101010101010101010110, 3'b000}); // 150: fn=  SUB, a=0x00000000, b=0xaaaaaaaa, y=0x55555556
	test_case({6'b010001, 32'b00000000000000000000000000000000, 32'b01010101010101010101010101010101}, {32'b10101010101010101010101010101011, 3'b001}); // 151: fn=  SUB, a=0x00000000, b=0x55555555, y=0xaaaaaaab
	test_case({6'b010001, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000001, 3'b000}); // 152: fn=  SUB, a=0x00000001, b=0x00000000, y=0x00000001
	test_case({6'b010001, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000000, 3'b100}); // 153: fn=  SUB, a=0x00000001, b=0x00000001, y=0x00000000
	test_case({6'b010001, 32'b00000000000000000000000000000001, 32'b11111111111111111111111111111111}, {32'b00000000000000000000000000000010, 3'b000}); // 154: fn=  SUB, a=0x00000001, b=0x-0000001, y=0x00000002
	test_case({6'b010001, 32'b00000000000000000000000000000001, 32'b10101010101010101010101010101010}, {32'b01010101010101010101010101010111, 3'b000}); // 155: fn=  SUB, a=0x00000001, b=0xaaaaaaaa, y=0x55555557
	test_case({6'b010001, 32'b00000000000000000000000000000001, 32'b01010101010101010101010101010101}, {32'b10101010101010101010101010101100, 3'b001}); // 156: fn=  SUB, a=0x00000001, b=0x55555555, y=0xaaaaaaac
	test_case({6'b010001, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000000}, {32'b11111111111111111111111111111111, 3'b001}); // 157: fn=  SUB, a=0x-0000001, b=0x00000000, y=0xffffffff
	test_case({6'b010001, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000001}, {32'b11111111111111111111111111111110, 3'b001}); // 158: fn=  SUB, a=0x-0000001, b=0x00000001, y=0xfffffffe
	test_case({6'b010001, 32'b11111111111111111111111111111111, 32'b11111111111111111111111111111111}, {32'b00000000000000000000000000000000, 3'b100}); // 159: fn=  SUB, a=0x-0000001, b=0x-0000001, y=0x00000000
	test_case({6'b010001, 32'b11111111111111111111111111111111, 32'b10101010101010101010101010101010}, {32'b01010101010101010101010101010101, 3'b000}); // 160: fn=  SUB, a=0x-0000001, b=0xaaaaaaaa, y=0x55555555
	test_case({6'b010001, 32'b11111111111111111111111111111111, 32'b01010101010101010101010101010101}, {32'b10101010101010101010101010101010, 3'b001}); // 161: fn=  SUB, a=0x-0000001, b=0x55555555, y=0xaaaaaaaa
	test_case({6'b010001, 32'b10101010101010101010101010101010, 32'b00000000000000000000000000000000}, {32'b10101010101010101010101010101010, 3'b001}); // 162: fn=  SUB, a=0xaaaaaaaa, b=0x00000000, y=0xaaaaaaaa
	test_case({6'b010001, 32'b10101010101010101010101010101010, 32'b00000000000000000000000000000001}, {32'b10101010101010101010101010101001, 3'b001}); // 163: fn=  SUB, a=0xaaaaaaaa, b=0x00000001, y=0xaaaaaaa9
	test_case({6'b010001, 32'b10101010101010101010101010101010, 32'b11111111111111111111111111111111}, {32'b10101010101010101010101010101011, 3'b001}); // 164: fn=  SUB, a=0xaaaaaaaa, b=0x-0000001, y=0xaaaaaaab
	test_case({6'b010001, 32'b10101010101010101010101010101010, 32'b10101010101010101010101010101010}, {32'b00000000000000000000000000000000, 3'b100}); // 165: fn=  SUB, a=0xaaaaaaaa, b=0xaaaaaaaa, y=0x00000000
	test_case({6'b010001, 32'b10101010101010101010101010101010, 32'b01010101010101010101010101010101}, {32'b01010101010101010101010101010101, 3'b010}); // 166: fn=  SUB, a=0xaaaaaaaa, b=0x55555555, y=0x55555555
	test_case({6'b010001, 32'b01010101010101010101010101010101, 32'b00000000000000000000000000000000}, {32'b01010101010101010101010101010101, 3'b000}); // 167: fn=  SUB, a=0x55555555, b=0x00000000, y=0x55555555
	test_case({6'b010001, 32'b01010101010101010101010101010101, 32'b00000000000000000000000000000001}, {32'b01010101010101010101010101010100, 3'b000}); // 168: fn=  SUB, a=0x55555555, b=0x00000001, y=0x55555554
	test_case({6'b010001, 32'b01010101010101010101010101010101, 32'b11111111111111111111111111111111}, {32'b01010101010101010101010101010110, 3'b000}); // 169: fn=  SUB, a=0x55555555, b=0x-0000001, y=0x55555556
	test_case({6'b010001, 32'b01010101010101010101010101010101, 32'b10101010101010101010101010101010}, {32'b10101010101010101010101010101011, 3'b011}); // 170: fn=  SUB, a=0x55555555, b=0xaaaaaaaa, y=0xaaaaaaab
	test_case({6'b010001, 32'b01010101010101010101010101010101, 32'b01010101010101010101010101010101}, {32'b00000000000000000000000000000000, 3'b100}); // 171: fn=  SUB, a=0x55555555, b=0x55555555, y=0x00000000
	test_case({6'b000011, 32'b00000000000000000000000000000101, 32'b11011110101011011011111011101111}, {32'b00000000000000000000000000000000, 3'b000}); // 172: fn=CMPEQ, a=0x00000005, b=0xdeadbeef, y=0x00000000
	test_case({6'b000101, 32'b00000000000000000000000000000101, 32'b11011110101011011011111011101111}, {32'b00000000000000000000000000000000, 3'b000}); // 173: fn=CMPLT, a=0x00000005, b=0xdeadbeef, y=0x00000000
	test_case({6'b000111, 32'b00000000000000000000000000000101, 32'b11011110101011011011111011101111}, {32'b00000000000000000000000000000000, 3'b000}); // 174: fn=CMPLE, a=0x00000005, b=0xdeadbeef, y=0x00000000
	test_case({6'b000011, 32'b00010010001101000101011001111000, 32'b00010010001101000101011001111000}, {32'b00000000000000000000000000000001, 3'b100}); // 175: fn=CMPEQ, a=0x12345678, b=0x12345678, y=0x00000001
	test_case({6'b000101, 32'b00010010001101000101011001111000, 32'b00010010001101000101011001111000}, {32'b00000000000000000000000000000000, 3'b100}); // 176: fn=CMPLT, a=0x12345678, b=0x12345678, y=0x00000000
	test_case({6'b000111, 32'b00010010001101000101011001111000, 32'b00010010001101000101011001111000}, {32'b00000000000000000000000000000001, 3'b100}); // 177: fn=CMPLE, a=0x12345678, b=0x12345678, y=0x00000001
	test_case({6'b000011, 32'b10000000000000000000000000000000, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000000, 3'b010}); // 178: fn=CMPEQ, a=0x80000000, b=0x00000001, y=0x00000000
	test_case({6'b000101, 32'b10000000000000000000000000000000, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000001, 3'b010}); // 179: fn=CMPLT, a=0x80000000, b=0x00000001, y=0x00000001
	test_case({6'b000111, 32'b10000000000000000000000000000000, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000001, 3'b010}); // 180: fn=CMPLE, a=0x80000000, b=0x00000001, y=0x00000001
	test_case({6'b000011, 32'b11011110101011011011111011101111, 32'b00000000000000000000000000000101}, {32'b00000000000000000000000000000000, 3'b001}); // 181: fn=CMPEQ, a=0xdeadbeef, b=0x00000005, y=0x00000000
	test_case({6'b000101, 32'b11011110101011011011111011101111, 32'b00000000000000000000000000000101}, {32'b00000000000000000000000000000001, 3'b001}); // 182: fn=CMPLT, a=0xdeadbeef, b=0x00000005, y=0x00000001
	test_case({6'b000111, 32'b11011110101011011011111011101111, 32'b00000000000000000000000000000101}, {32'b00000000000000000000000000000001, 3'b001}); // 183: fn=CMPLE, a=0xdeadbeef, b=0x00000005, y=0x00000001
	test_case({6'b000011, 32'b01111111111111111111111111111111, 32'b11111111111111111111111111111111}, {32'b00000000000000000000000000000000, 3'b011}); // 184: fn=CMPEQ, a=0x7fffffff, b=0xffffffff, y=0x00000000
	test_case({6'b000101, 32'b01111111111111111111111111111111, 32'b11111111111111111111111111111111}, {32'b00000000000000000000000000000000, 3'b011}); // 185: fn=CMPLT, a=0x7fffffff, b=0xffffffff, y=0x00000000
	test_case({6'b000111, 32'b01111111111111111111111111111111, 32'b11111111111111111111111111111111}, {32'b00000000000000000000000000000000, 3'b011}); // 186: fn=CMPLE, a=0x7fffffff, b=0xffffffff, y=0x00000000
	$display("");
    $finish;
end


beta_alu dut (
	.a(a),
	.b(b),
    .fn(fn),
    .y(y)
);

endmodule
